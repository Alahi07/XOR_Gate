// Code your design here
module xorgate(
  input a,b,
  output y);
  assign y= a^b;
endmodule


